`include "verif.svh"


`define clk tb.clock
`define rst tb.reset